-- ------------------------------------------------------------------
-- --  _____       ______  _____                                   --
-- -- |_   _|     |  ____|/ ____|                                  --
-- --   | |  _ __ | |__  | (___    Institute of Embedded Systems   --
-- --   | | | '_ \|  __|  \___ \   Zurich University of            --
-- --  _| |_| | | | |____ ____) |  Applied Sciences                --
-- -- |_____|_| |_|______|_____/   8401 Winterthur, Switzerland    --
-- ------------------------------------------------------------------
--! @file crc5_gen.vhd
--! @author scso <scso@zhaw.ch>
--! @copyright 2022 ZHAW Institute of Embedded Systems
--! @date 2022-05-06
--! @brief generates 5 bit crc for up to 4 bytes of data using a lut generated by the 0x2b polynom
--! polynom has been taken from https://users.ece.cmu.edu/~koopman/crc/hd4.html
--! 
---------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Entity Declaration 
-------------------------------------------
entity crc5_gen is
    port (
        clk      : in  std_logic;
        rst_n    : in  std_logic;
        enable_i : in  std_logic; -- triggeres a crc 
        clear_i  : in  std_logic; -- clears the cached crc value
        crc_i    : in  std_logic; -- signals whether the data_i hold an already generated crc that should be used for validation
        data_i   : in  std_logic_vector(7 downto 0);
        crc_o    : out std_logic_vector(4 downto 0)
    );
end crc5_gen;

-- Architecture Declaration
-------------------------------------------
architecture rtl of crc5_gen is
    -- Component Declarations
    -------------------------------------------

    -- Signals & Constants Declaration
    -------------------------------------------
    type vec_arr_t is array (0 to 255) of std_logic_vector(7 downto 0);


    constant lut_crc5 : vec_arr_t := (
        x"00", x"0b", x"16", x"1d", x"07", x"0c", x"11", x"1a", x"0e", x"05",
        x"18", x"13", x"09", x"02", x"1f", x"14", x"1c", x"17", x"0a", x"01",
        x"1b", x"10", x"0d", x"06", x"12", x"19", x"04", x"0f", x"15", x"1e",
        x"03", x"08", x"13", x"18", x"05", x"0e", x"14", x"1f", x"02", x"09",
        x"1d", x"16", x"0b", x"00", x"1a", x"11", x"0c", x"07", x"0f", x"04",
        x"19", x"12", x"08", x"03", x"1e", x"15", x"01", x"0a", x"17", x"1c",
        x"06", x"0d", x"10", x"1b", x"0d", x"06", x"1b", x"10", x"0a", x"01",
        x"1c", x"17", x"03", x"08", x"15", x"1e", x"04", x"0f", x"12", x"19",
        x"11", x"1a", x"07", x"0c", x"16", x"1d", x"00", x"0b", x"1f", x"14",
        x"09", x"02", x"18", x"13", x"0e", x"05", x"1e", x"15", x"08", x"03",
        x"19", x"12", x"0f", x"04", x"10", x"1b", x"06", x"0d", x"17", x"1c",
        x"01", x"0a", x"02", x"09", x"14", x"1f", x"05", x"0e", x"13", x"18",
        x"0c", x"07", x"1a", x"11", x"0b", x"00", x"1d", x"16", x"1a", x"11",
        x"0c", x"07", x"1d", x"16", x"0b", x"00", x"14", x"1f", x"02", x"09",
        x"13", x"18", x"05", x"0e", x"06", x"0d", x"10", x"1b", x"01", x"0a",
        x"17", x"1c", x"08", x"03", x"1e", x"15", x"0f", x"04", x"19", x"12",
        x"09", x"02", x"1f", x"14", x"0e", x"05", x"18", x"13", x"07", x"0c",
        x"11", x"1a", x"00", x"0b", x"16", x"1d", x"15", x"1e", x"03", x"08",
        x"12", x"19", x"04", x"0f", x"1b", x"10", x"0d", x"06", x"1c", x"17",
        x"0a", x"01", x"17", x"1c", x"01", x"0a", x"10", x"1b", x"06", x"0d",
        x"19", x"12", x"0f", x"04", x"1e", x"15", x"08", x"03", x"0b", x"00",
        x"1d", x"16", x"0c", x"07", x"1a", x"11", x"05", x"0e", x"13", x"18",
        x"02", x"09", x"14", x"1f", x"04", x"0f", x"12", x"19", x"03", x"08",
        x"15", x"1e", x"0a", x"01", x"1c", x"17", x"0d", x"06", x"1b", x"10",
        x"18", x"13", x"0e", x"05", x"1f", x"14", x"09", x"02", x"16", x"1d",
        x"00", x"0b", x"11", x"1a", x"07", x"0c");
    signal crc : std_logic_vector(7 downto 0) := (others => '0');
-- Begin Architecture
-------------------------------------------
begin
    --------------------------------------------------
    -- PROCESS FOR REGISTERS
    --------------------------------------------------
    clocking : process (clk, rst_n)
        variable v_data : std_logic_vector(data_i'range) := (others => '0');
    begin
        if rst_n = '0' then
            crc <= (others => '0');
        elsif rising_edge(clk) then
            if enable_i = '1' then
                if crc_i = '1' then
                    -- if crc is enterd for crc validation, it is only 6 bit long and needs to be MSB aligned
                    v_data := data_i(4 downto 0)&"000";
                else 
                    v_data := data_i;
                end if;

                if clear_i = '1' then
                    crc <= lut_crc5(to_integer(unsigned(v_data xor x"00")));
                else
                    -- discard MSB of cached crc and pad with LSB 0
                    crc <= lut_crc5(to_integer(unsigned(v_data xor crc(4 downto 0)&"000")));
                end if;
            elsif clear_i = '1' then
                crc <= x"00";
            end if;
        end if;
    end process clocking;

    --------------------------------------------------
    -- CONCURRENT ASSIGNMENTS
    --------------------------------------------------
    crc_o <= crc(4 downto 0);
------------------------------------------- 
-- End Architecture 
------------------------------------------- 
end rtl;
